module()


endmodule
