module()
input a;

endmodule
